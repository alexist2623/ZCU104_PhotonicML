{
    "verilog" : {
        "name" : "HDMIController",
        "top": "HDMIController.sv",
        "files" : [
            "HDMIController/HDMIController.sv"
        ]
    }
}